module instruction_memory(input logic[7:0] PC,
                        output logic[23:0] Instr);
