`timescale 1ps/1ps
`include "pc.sv"
